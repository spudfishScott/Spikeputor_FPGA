-- megafunction wizard: %RAM: 1-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altsyncram 

-- ============================================================
-- File Name: RAM.vhd
-- Megafunction Name(s):
--          altsyncram
--
-- Simulation Library Files(s):
--          altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.1.0 Build 162 10/23/2013 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


-- RAM module - outputs words of 16 bits each - single port, NUM_WORDS must be powers of 2
LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY RAM IS
    GENERIC (
        NUM_WORDS  : INTEGER := 16384;          -- 32K bytes = 16K words of 16 bits each
        ADDR_WIDTH : INTEGER := 14              -- 14 bits to address 16K words
    );

    PORT (
        clock       : IN STD_LOGIC  := '1';

        address     : IN STD_LOGIC_VECTOR (ADDR_WIDTH-1 DOWNTO 0);
        data        : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        wren        : IN STD_LOGIC  := '0';

        q           : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
    );
END RAM;

ARCHITECTURE SYN OF RAM IS
    SIGNAL sub_wire0    : STD_LOGIC_VECTOR (15 DOWNTO 0);                   -- output is latched

BEGIN
    q    <= sub_wire0(15 DOWNTO 0);

    altsyncram_component : altsyncram
    GENERIC MAP (
        clock_enable_input_a => "BYPASS",
        clock_enable_output_a => "BYPASS",
        intended_device_family => "Cyclone III",
        lpm_hint => "ENABLE_RUNTIME_MOD=NO",
        lpm_type => "altsyncram",
        numwords_a => NUM_WORDS,
        operation_mode => "SINGLE_PORT",
        outdata_aclr_a => "NONE",
        outdata_reg_a => "CLOCK0",
        power_up_uninitialized => "FALSE",
        read_during_write_mode_port_a => "NEW_DATA_NO_NBE_READ",
        widthad_a => ADDR_WIDTH,
        width_a => 16,
        width_byteena_a => 1
    )
    PORT MAP (
        address_a => address,
        clock0 => clock,
        data_a => data,
        wren_a => wren,
        q_a => sub_wire0
    );

END SYN;
