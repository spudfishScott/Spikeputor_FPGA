-- Spikeputor Control Logic and Memory Wishbone Interface Master
-- Data and ADDRESS buses are 16 bits wide
-- Each CPU instruction cycle can be up to three read/writes, so execute them in a single wishbone BLOCK READ/WRITE cycle
-- ACK_I is the only termination signal currently supported. RTY_I and ERR_I are not supported.

-- Contains the INST, CONST, and PC registers
-- Also contains the state machine for fetching instructions and constants from memory
-- and executing instructions, including memory read and write operations.
-- Uses a simple 4-state FSM to manage instruction fetch, constant fetch, and execution phases (with out without memory r/w command)
-- Includes a PHASE output to indicate current phase of instruction cycle for display purposes
-- Memory interface is a Wishbone Master interface
-- Inputs from ALU and Register File, outputs to Register File and ALU control signals
-- Memory write data is directly from Register File Channel B output (MWDATA)
-- Memory Read Data is output to MRDATA signal
-- Program Counter (PC) is incremented by 2 for each instruction, unless a branch or jump occurs
-- On reset, PC is set to the RESET_VECTOR address (xF000)
-- Instruction format:
--     Bits 15-11: ALU Opcode
--     Bit 10:    '1' if instruction has a constant (CONST), '0' if no constant
--     Bit 9:     '1' if instruction is a memory (LD, LDR, ST) or branch (JMP, BEQ, BNE) operation, '0' for other instructions
--     Bits 8-6:  Register Operand B or Memory/Branch opcode
--                For memory operations:
--                  "010" for LD and LDC instructions
--                  "110" for LDR instruction
--                  "011" for ST and STC instructions
--                For branch instructions:
--                  "000" = JMP (unconditional)
--                  "100" = BEQ (branch if zero)
--                  "101" = BNE (branch if not zero)
--     Bits 5-3:  Register Operand C
--     Bits 2-0:  Register Operand A - directly to Channel A of Register File
-- ALU Control signals:
    -- ALUFN: INST(15 downto 11)
    -- ASEL:  INST(8) AND INST(9)
    -- BSEL:  INST(10)
-- Register File Control signals:
    -- WERF:  '1' to write to register file, '0' otherwise
    -- RBSEL: '0' to select OPB, '1' to select OPC for Channel B output
    -- WDSEL: "01" to select ALU output, "00" to select PC+2, "10" to select Memory Read Data
    -- OPA:   INST(2 downto 0)
    -- OPB:   INST(8 downto 6)
    -- OPC:   INST(5 downto 3)

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Types.all;

entity CTRL_WSH_M is
    port (
        -- SYSCON inputs
        CLK         : in std_logic;
        RST_I       : in std_logic;

        -- Wishbone signals for memory interface
        -- handshaking signals
        WBS_CYC_O   : out std_logic;
        WBS_STB_O   : out std_logic;
        WBS_ACK_I   : in std_logic;

        -- memory read/write signals
        WBS_ADDR_O  : out std_logic_vector(15 downto 0);    -- lsb is ignored, but it is still part of the address bus
        WBS_DATA_O  : out std_logic_vector(15 downto 0);    -- data output to provider
        WBS_DATA_I  : in std_logic_vector(15 downto 0);     -- data input from provider
        WBS_WE_O    : out std_logic;                        -- write enable output - write when high, read when low

        -- Spikeputor Signals
            -- Data outputs from Control Logic to other modules
        INST    : out std_logic_vector(15 downto 0);                      -- instruction fetched from memory - for display only
        CONST   : out std_logic_vector(15 downto 0);                      -- constant fetched from memory
        PC      : out std_logic_vector(15 downto 0);                      -- program counter
        PC_INC  : out std_logic_vector(15 downto 0);                      -- incremented program counter
        MRDATA  : out std_logic_vector(15 downto 0);                      -- memory read data

            -- Control signals from Control Logic to RegFile
        WERF    : out std_logic;                                          -- Write Enable Register File - '1' to write to register file
        RBSEL   : out std_logic;                                          -- Register Channel B Select - '0' for OPB, '1' for OPC
        WDSEL   : out std_logic_vector(1 downto 0);                       -- Write Data Select - "01" for ALU, "00" for PC+2, "10" for Memory Read Data
        OPA     : out std_logic_vector(2 downto 0);                       -- Register Operand A
        OPB     : out std_logic_vector(2 downto 0);                       -- Register Operand B
        OPC     : out std_logic_vector(2 downto 0);                       -- Register Operand C

            -- Control signals from Control Logic to ALU
        ALUFN   : out std_logic_vector(4 downto 0);                       -- ALU Function select - opcode from instruction
        ASEL    : out std_logic;                                          -- ALU A input select - '0' for REGFile Channel A, '1' for PC+2
        BSEL    : out std_logic;                                          -- ALU B input select - '0' for REGFile Channel B, '1' for CONST

            -- Inputs to Control Logic from other modules
        ALU_OUT : in std_logic_vector(15 downto 0);                       -- ALU output
        MWDATA  : in std_logic_vector(15 downto 0);                       -- memory write data - Register Channel B output
        Z       : in std_logic;                                           -- Zero flag from RegFile Channel A

        PHASE   : out std_logic_vector(1 downto 0)                        -- current phase of instruction cycle
    );
end CTRL_WSH_M;

architecture rtl of CTRL_WSH_M is

    -- internal signals
    constant RESET_VECTOR : std_logic_vector(15 downto 0) := x"F000";   -- reset vector address

    -- internal registers to hold outputs
    signal INST_reg    : std_logic_vector(15 downto 0) := (others => '0');   -- instruction fetched from memory
    signal CONST_reg   : std_logic_vector(15 downto 0) := (others => '0');   -- constant fetched from memory
    signal PC_reg      : std_logic_vector(15 downto 0) := (others => '0');   -- program counter
    signal PC_INC_calc : std_logic_vector(15 downto 0) := (others => '0');   -- incremented program counter
    signal MRDATA_reg  : std_logic_vector(15 downto 0) := (others => '0');   -- memory read data
    
    signal RBSEL_sig   : std_logic := '0';                                   -- Register Channel B Select - '0' for OPB, '1' for OPC
    signal WERF_sig    : std_logic := '0';                                   -- Write Enable for Register File - on during execute phase if instruction is not a store (ST command)
    signal WDSEL_sig   : std_logic_vector(1 downto 0) := (others => '0');    -- Write Data Select - "01" for ALU, "00" for PC+2, "10" for Memory Read Data
    signal OPA_sig     : std_logic_vector(2 downto 0) := (others => '0');    -- Register Operand A
    signal OPB_sig     : std_logic_vector(2 downto 0) := (others => '0');    -- Register Operand B
    signal OPC_sig     : std_logic_vector(2 downto 0) := (others => '0');    -- Register Operand C

    signal ALUFN_sig   : std_logic_vector(4 downto 0) := (others => '0');    -- ALU Function select - opcode from instruction
    signal ASEL_sig    : std_logic := '0';                                   -- ALU A input select - '0' for REGFile Channel A, '1' for PC+2
    signal BSEL_sig    : std_logic := '0';                                   -- ALU B input select - '0' for REGFile Channel B, '1' for CONST

    -- state machine
    type fsm_main is (ST_FETCH_I, ST_FETCH_C, ST_EXECUTE, ST_EXECUTE_RW);
    signal st_main : fsm_main := ST_FETCH_I;

begin
    -- Spikeputor control outputs, including control signals for ALU and Register File
    PC          <= PC_reg;                                                  -- program counter
    PC_INC      <= PC_INC_calc;                                             -- incremented program counter
    INST        <= INST_reg;                                                -- instruction fetched from memory
    CONST       <= CONST_reg;                                               -- constant fetched from memory
    MRDATA      <= MRDATA_reg;                                              -- memory read data
    RBSEL       <= RBSEL_sig;                                               -- Register Channel B Select - '0' for OPB, '1' for OPC
    WERF        <= WERF_sig;                                                -- Write Enable for Register File - on during execute phase if instruction is not a store (ST command)
    WDSEL       <= WDSEL_sig;                                               -- Write Data Select - "01" for ALU, "00" for PC+2, "10" for Memory Read Data
    OPA         <= OPA_sig;                                                 -- Register Operand A
    OPB         <= OPB_sig;                                                 -- Register Operand B
    OPC         <= OPC_sig;                                                 -- Register Operand C
    ALUFN       <= ALUFN_sig;                                               -- ALU Function select - opcode from instruction
    ASEL        <= ASEL_sig;                                                -- ALU A input select - '0' for REGFile Channel A, '1' for PC+2
    BSEL        <= BSEL_sig;                                                -- ALU B input select - '0' for REGFile Channel B

    PHASE       <=  "00" when st_main = ST_FETCH_I else                     -- current phase of instruction cycle for display purposes
                    "01" when st_main = ST_FETCH_C else
                    "10" when st_main = ST_EXECUTE else
                    "11" when st_main = ST_EXECUTE_RW else
                    "00";  -- should never occur, default to fetch instruction phase

    PC_INC_calc <= std_logic_vector(unsigned(PC_reg) + 2);

    process(clk)
    begin
        if rising_edge(clk) then
            if RST_I = '1' then
                -- reset state
                st_main <= ST_FETCH_I;          -- start by fetching instruction
                PC_reg <= RESET_VECTOR;         -- set PC to reset vector

                 -- clear wishbone signals
                WBS_CYC_O <= '0';               -- clear wishbone handshake signals
                WBS_STB_O <= '0';
                WBS_WE_O <= '0';
                WBS_ADDR_O <= RESET_VECTOR;     -- set address to reset vector
                WBS_DATA_O <= (others => '0');  -- clear data output
            else
                -- normal operation
                WBS_DATA_O <= MWDATA;           -- data output is directly from Register File Channel B output when reset = '0'
                WERF_sig <= '0';                -- clear write enable signal until we reach execute state

                case st_main is
                    when ST_FETCH_I =>
                        -- fetch instruction from memory at address PC
                        WBS_ADDR_O <= PC_reg;           -- set address to PC
                        WBS_CYC_O <= '1';               -- initiate wishbone cycle
                        WBS_STB_O <= '1';               -- strobe to indicate valid address and start memory read
                        WBS_WE_O <= '0';                -- read operation
                        if WBS_ACK_I = '1' then     -- wait for acknowledge from memory
                            INST_reg <= WBS_DATA_I;     -- latch instruction
                            -- decode instruction to set control signals for ALU and Register File
                            ALUFN_sig <= WBS_DATA_I(15 downto 11);
                            ASEL_sig <= WBS_DATA_I(8) AND WBS_DATA_I(9);  -- ASEL = 1 for PC+2 (for memory and branching instructions), else 0 for RegFile Channel A
                            BSEL_sig <= WBS_DATA_I(10);                   -- BSEL = 1 for CONST (for instructions that get a constant), else 0 for RegFile Channel B
                            OPA_sig <= WBS_DATA_I(2 downto 0);            -- OPA is always bits 2-0
                            OPB_sig <= WBS_DATA_I(8 downto 6);            -- OPB is always bits 8-6
                            OPC_sig <= WBS_DATA_I(5 downto 3);            -- OPC is always bits 5-3
                            
                            if WBS_DATA_I(8 downto 6) = "011" then        -- if ST instruction, select OPC for RegFile Channel B output
                                RBSEL_sig <= '1';
                            else
                                RBSEL_sig <= '0';
                            end if;

                            WBS_STB_O <= '0';           -- deassert strobe - end read phase
                            if WBS_DATA_I(10) = '1' then    -- instruction bit 10 indicates if there is a constant to fetch
                                st_main <= ST_FETCH_C;          -- instruction has constant
                                PC_reg <= PC_INC_calc;          -- increment PC for constant
                            else
                                PC_reg <= PC_reg;
                                st_main <= ST_EXECUTE;          -- no constant, execute directly (keeping PC unchanged)
                            end if;
                        else                        -- stall until ack received
                            st_main <= ST_FETCH_I;
                        end if;

                    when ST_FETCH_C =>
                        -- fetch constant from memory at now incremented PC
                        WBS_ADDR_O <= PC_reg;           -- set address to PC
                        WBS_STB_O <= '1';               -- strobe to indicate valid address and start memory read
                        WBS_WE_O <= '0';                -- read operation
                        if WBS_ACK_I = '1' then
                            CONST_reg <= WBS_DATA_I;    -- latch constant
                            WBS_STB_O <= '0';           -- deassert strobe - end read phase
                            st_main <= ST_EXECUTE;      -- proceed to execute instruction
                        else
                            st_main <= ST_FETCH_C;  -- stall until ack received
                        end if;

                    when ST_EXECUTE =>
                        -- execute instruction
                        WERF_sig <= NOT RBSEL_sig;                      -- set WERF flag on execute - write to register file if not a store (ST command)
                                                                        -- set WDSEL
                        if (INST_reg(9) = '1' AND INST_reg(7 downto 6) = "10") then
                            WDSEL_sig <= "10";                         -- use Memory Read Data as Register Input for LD and LDR instructions
                        elsif (INST_reg(9) = '1' AND INST_reg(7) = '0') then
                            WDSEL_sig <= "00";                         -- use PC+2 as Register Input for Branch Instructions
                        else
                            WDSEL_sig <= "01";                         -- use ALU Output as Register Input for all other instructions
                        end if;

                        if (INST_reg(9) AND INST_reg(7)) = '1' then     -- operation requires memory read or write (LD, LDR, or ST - formerly MASEL = 1)
                            WBS_ADDR_O <= ALU_OUT;                          -- address is ALU output
                            WBS_STB_O <= '1';                               -- strobe to indicate valid address and start memory read/write
                            if (INST_reg(9) AND RBSEL_sig) = '1' then       -- write to memory on ST command (formerly MWR = 1), otherwise read
                                WBS_WE_O <= '1';
                            else
                                WBS_WE_O <= '0';
                            end if;
                            st_main <= ST_EXECUTE_RW;       -- wait in execute_rw state until ack received
                        else                            -- other instructions - do not need to read or write to memory
                            if ((INST_reg(9) = '1') AND                   -- check to see if the branch should be taken (formerly JT = 1)
                                    ((INST_reg(8 downto 6) = "000") OR                        -- unconditional jump (JMP)
                                    (INST_reg(8 downto 6) = "100" AND Z_sig = '1') OR         -- branch if equal to zero (BEQ)
                                    (INST_reg(8 downto 6) = "101" AND Z_sig = '0'))) then     -- branch if not equal to zero (BNE)
                                        PC_reg <= ALU_OUT;          -- set PC to address in ALU output to jump
                            else
                                        PC_reg <= PC_INC_calc;      -- increment PC by 2 for next instruction
                            end if;
                            WBS_CYC_O <= '0';               -- end wishbone cycle
                            st_main <= ST_FETCH_I;          -- go back to fetch next instruction, no wishbone cycle needed
                        end if;

                    when ST_EXECUTE_RW =>
                        -- wait state for memory read or write operation to complete
                        if WBS_ACK_I = '1' then         -- wait for acknowledge from memory and handle read or write completion
                            if (INST_reg(9) AND RBSEL_sig) = '0' then   -- if not a store command (formerly MRW = 0), it is a memory read operation
                                MRDATA_reg <= WBS_DATA_I;   -- latch memory read data for read operation
                            else 
                                WBS_WE_O <= '0';            -- deassert write enable after write operation
                            end if;

                            PC_reg <= PC_INC_calc;      -- increment PC by 2 for next instruction
                            WBS_STB_O <= '0';           -- deassert strobe
                            WBS_CYC_O <= '0';           -- end wishbone cycle
                            st_main <= ST_FETCH_I;      -- go back to fetch next instruction
                        else
                            st_main <= ST_EXECUTE_RW;   -- stall until ack received
                        end if;

                    when others =>                  -- should never occur
                        st_main <= ST_FETCH_I;          -- default to fetch instruction state
                end case;
            end if;
        end if;
    end process;

end rtl;