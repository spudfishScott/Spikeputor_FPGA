-- This is a Wishbone address comparitor to route bus inputs to a variety of provider models
-- Inputs are:
--  TGA_I  - from the master arbiter (either extended address via SEGMENT register or 0)
--  ADDR_I - from the master arbiter
--  WE_I   - from the master arbiter
--  STB_I  - from the master arbiter
--  TGD_I  - route the data bus to update the SEGMENT register
        --      If TGA_I is not 0, RAM?ROM is determined by msb (bit 23) of ADDR_I (1 = ROM, 0 = RAM)
--  Px_DATA_O - data output from each provider
--
-- In addition to standard RAM (P0), SDRAM (P10), and ROM (P1), the following providers are accessed through specific addresses, which override the above:
--  GPO (P2)        read/write location 0x7FFC
--  GPI (P3)        read only location 0x7FFE - writing goes nowhere
--  SOUND (P4)      read/write location 0x7FAC
--  VIDEO (P5)      read/write to video coprocessor - locations TBD
--  SERIAL (P6)     serial in/serial out - locations TBD
--  STORAGE (P7)    read/write to SD card filesystem - locations TBD (might be coupled to DMA)
--  KEYBOARD (P8)   read keyboard input buffer (maybe mouse one day as well)
--  SEGMENT (P9)    read/write to segment register, which might be used to expand the total amount of RAM available - locations TBD
--  MATH (P11)      floating point unit - locations TBD

-- Outputs are:
--  Individual provider select signals, which go to provider STB_I inputs
--  DATA_O - wired to all of the master DATA_I inputs

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Types.all;

entity WSH_ADDR is
    port (
        -- Wishbone Control Signals
        ADDR_I      : in std_logic_vector(23 downto 0);     -- standard address bus - bottom 16 bits is on Segment 0, msb = ROM/RAM for extended memory, bits 22->16 = segment number
        WE_I        : in std_logic;                         -- write enable flag
        STB_I       : in std_logic;                         -- wishbone strobe signal
        TGD_I       : in std_logic;                         -- when TGD_I and WE_I are high, route to P9, SEGMENT write

        -- Data out from providers
        P0_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from RAM (P0) 0x0000-0xDFFF
        P1_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from ROM (P1) 0xE000-0xFFFF, 0x810000-0xBFFFFF
        P2_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from GPO (P2)
        P3_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from GPI (P3)
        P4_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from SOUND (P4)
        P5_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from VIDEO (P5)
        P6_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from SERIAL (P6)
        P7_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from STORAGE (P7)
        P8_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from KEYBOARD (P8)
        P9_DATA_O   : in std_logic_vector(15 downto 0);     -- Data Output from SEGMENT (P9)
        P10_DATA_O  : in std_logic_vector(15 downto 0);     -- Data Output from SDRAM (P10) 0x010000-0x7FFFFF
        P11_DATA_O  : in std_logic_vector(15 downto 0);     -- Data Output from MATH (P11)

        -- Output signals
        DATA_O      : out std_logic_vector(15 downto 0);    -- Wishbone data bus output
        STB_SEL     : out std_logic_vector(11 downto 0)     -- One hot strobe selector for provider STB_I signals
    );
end WSH_ADDR;

architecture RTL of WSH_ADDR is
                            -- (map low byte of address to video coprocessor registers, except 0x00 => STATUS, and protect against registers that should not be exposed)
    constant VIDEO_ADDR     : std_logic_vector(15 downto 0) := x"FF00"; -- VIDEO address start (0xFF00-0xFFDF)
    constant KEYBOARD_ADDR  : std_logic_vector(15 downto 0) := x"FFF0"; -- keyboard address - read only
    constant GPO_ADDR       : std_logic_vector(15 downto 0) := x"FFF1"; -- GPO address - read/write
    constant GPI_ADDR       : std_logic_vector(15 downto 0) := x"FFF2"; -- GPI address - read only

-- math fpu - two 32-bit input addresses, one 32-bit output addresses, one control/status address - 7 total (0xFFE0-0xFFE6)
-- sound - use VGA output for sound? three voices, 4-bits each. So one address for volume and waveform control of all three voices, one address for frequency control for each voice - 4 total
-- serial - one address I/O
-- storage - one address I/O

    signal p_sel   : integer range 0 to 11 := 0;                        -- provider selector index
    signal ram_e   : std_logic := '0';                                  -- FPGA RAM selected
    signal spec    : std_logic := '0';                                  -- special location (p2-p9)
    signal sdram_e : std_logic := '0';                                  -- sdram selected
    signal seg     : std_logic_vector(6 downto 0) := (others => '0');   -- segment portion of the full address
    signal p_addr  : std_logic_vector(15 downto 0) := (others => '0');  -- primary address portion of the full address
    signal p_oh    : std_logic_vector(11 downto 0) := (others => '0');  -- provider one-hot vector

begin
    seg    <= ADDR_I(22 downto 16);   -- extract segment identifier from full address
    p_addr <= ADDR_I(15 downto 0);    -- extract primary address from full address

    spec    <= '1' when seg = "0000000" AND p_addr(15 downto 8) = x"FF"                     -- special I/O address
                   else '0';
    ram_e   <= '1' when (seg  = "0000000" AND ADDR_I(15 downto 13) /= "111")                -- standard RAM:0x0000-0xDFFF, Segment 0
                   else '0';
    sdram_e <= '1' when (seg /= "0000000" AND ADDR_I(23) = '0')                             -- SDRAM: not segment 0 and not a ROM address
                   else '0';

    -- assign p_sel based on addressing logic described above
    p_sel <=    9 when TGD_I = '1' AND WE_I = '1'                                         -- write to SEGMENT when TDG and WE are set, pre-empts all other
        else    0 when ram_e = '1'                                                        -- standard RAM
        else    1 when spec = '0' AND ram_e = '0' AND sdram_e = '0'                       -- ROM if not a special I/O location and not a RAM location (including 0xE000-0xFFFF)
        else    2 when spec = '1' AND p_addr = GPO_ADDR                                   -- read/write GPO
        else    3 when spec = '1' AND p_addr = GPI_ADDR                                   -- read only GPI
        -- to do the rest 4, 6, 7, 11
        else    8 when spec = '1' AND p_addr = KEYBOARD_ADDR                              -- read only KEYBOARD
        else    5 when spec = '1' AND p_addr(15 downto 8) = VIDEO_ADDR(15 downto 8) 
                                  AND p_addr(7 downto 4) < x"E"                           -- VIDEO coprocessor if address matches video range (0xFF00 - 0xFFDF)
        else   10 when ram_e = '1'                                                        -- SDRAM when ram_e is '1' and we get here (segment /= 0 and not ROM or special)
        else    1;                                                                        -- default to read ROM

    -- output the correct data based on p_sel
    with (p_sel) select
        DATA_O <=
            P0_DATA_O  when 0,      -- RAM
            P1_DATA_O  when 1,      -- ROM
            P2_DATA_O  when 2,      -- GPO (including VFD text output?)
            P3_DATA_O  when 3,      -- GPI
            P4_DATA_O  when 4,      -- SOUND
            P5_DATA_O  when 5,      -- VIDEO
            P6_DATA_O  when 6,      -- SERIAL
            P7_DATA_O  when 7,      -- DISK STORAGE
            P8_DATA_O  when 8,      -- KEYBOARD
            P9_DATA_O  when 9,      -- SEGMENT
            P10_DATA_O when 10,     -- SDRAM
            P11_DATA_O when 11,     -- MATH FPU
            (others => '0') when others;

    -- Generate one-hot strobe signals for each provider based on p_sel
    with (p_sel) select
        p_oh <=
            "000000000001" when 0,
            "000000000010" when 1,
            "000000000100" when 2,
            "000000001000" when 3,
            "000000010000" when 4,
            "000000100000" when 5,
            "000001000000" when 6,
            "000010000000" when 7,
            "000100000000" when 8,
            "001000000000" when 9,
            "010000000000" when 10,
            "100000000000" when 11,
            "000000000000" when others;

    -- ouput STB_SEL based on the one-hot result and STB_I
    STB_SEL <= p_oh when STB_I = '1' else "000000000000";

end RTL;
