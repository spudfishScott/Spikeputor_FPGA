-- External interface to the Spiekputor DMA - mediated through a serial connection to the outside world
-- Sends external signals:
    -- Start (begin the DMA transaction)
    -- Write/nRead (1 = write, 0 = read)
    -- Start Address (Full 24 Bit: msb = ROM/RAM for extended memory, bits 22->16 = segment number , bits 15->0 = address)
    -- Length - Number of bytes to read - 16 bits
    -- Write Data  - 16 bits sent to Spikeputor memory
    -- Read Data - 16 bits sent from Spikeputor memory
    -- Write Ready - ready to send the next word to the Spikeputor
    -- Read Ready - ready to send the next word from the Spikeputor

-- External Interface sends Start signal when Write/Read, Start Address, and Length are valid
-- If read, DMA gets first word, sets DATA_OUT, strobes READY_OUT, External Interface behaves as below
-- If write, External Interface gets first word, sets WR_DATA strobes WR_READY, DMA behaves as below
-- Data transfer continues:
    -- For Read: 
        -- External Interface waits for RD_READY, then latches RD_DATA, sends out word through serial port, strobes WR_READY, then loops until LENGTH bytes have been recieved
        -- DMA reads memory, sets RD_DATA, waits for WR_READY, strobes RD_READY, then loops until LENGTH bytes have been sent
    -- For Write:
        -- External Interface gets next word of data, sets WR_DATA, waits for RD_READY, strobes WR_READY, then loops until LENGTH bytes have been sent
        -- DMA waits for WR_READY, then latches WR_DATA, writes it to Spikeputor, strobes RD_READY, loops until LENGTH bytes have been received

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity dma_uart_ctrl is
    generic (
        CLK_FREQ   : Integer := 50_000_000;                     -- clock frequency - default = 50 MHz
    );
    port (
        CLK        : in  std_logic;
        RST        : in  std_logic;

        -- UART interface
        RX_SERIAL  : in std_logic;                              -- serial data input
        TX_SERIAL  : out std_logic;                             -- serial data output

        -- control signals (from UART interface)
        START       : out std_logic;                            -- strobe to begin DMA transaction
        WR_RD       : out std_logic;                            -- Write / nRead (1 = Write to Spikeputor, 0 - Read from Spikeputor)
        ADDRESS     : out std_logic_vector(23 downto 0);        -- Start address (full 24 bit)
        LENGTH      : out std_logic_vector(15 downto 0);        -- Length in bytes to read/write
        WR_DATA     : out std_logic_vector(15 downto 0);        -- Data to send to Spikeputor
        WR_READY    : out std_logic;                            -- Strobed when WR_DATA is valid
        RD_DATA     : in std_logic_vector(15 downto 0);         -- Data to send from the Spikeputor
        RD_READY    : in std_logic;                             -- Strobed when RD_DATA is valid
        RESET_REQ   : out std_logic;                            -- Request to reset the spikeputor
    );
end entity dma_uart_ctrl;

architecture behavioral of dma_uart_ctrl is

    signal uart_rx_data : std_logic_vector(7 downto 0);         -- Data received from UART
    signal uart_rx_rdy  : std_logic;                            -- Strobed when a byte is ready to be read from UART
    signal uart_tx_data : std_logic_vector(7 downto 0);         -- Data to send through UART
    signal uart_tx_load : std_logic;                            -- Strobe to load data into UART transmitter
    signal uart_tx_busy : std_logic;                            -- Indicates if UART transmitter is busy

    --  CONSTANTS
    constant C_READ  : std_logic_vector(7 downto 0) := x"3E";  -- '>' READ
    constant C_WRITE : std_logic_vector(7 downto 0) := x"3C";  -- '<' WRITE
    constant C_RESET : std_logic_vector(7 downto 0) := x"21";  -- '!' RESET
    constant C_ACK   : std_logic_vector(7 downto 0) := x"2A";  -- '*' ACK

    -- internal signals, including state machine
    -- include preliminary values for all to help with fitter getting stuck
    type proto_fsm is (
        WAIT_START, ACK_READ, ACK_WRITE, ACK_RESET,
        HDR_0, HDR_1, HDR_2, HDR_3, HDR_4,
        LOAD_L, LOAD_H, SEND_L, SEND_H,
        ACK_DONE
    );
    signal p_state     : proto_fsm := WAIT_START;                           -- start in WAIT_START state

    signal address     : std_logic_vector(23 downto 0) := (others => '0');  -- full 24 bit address
    signal write_len   : unsigned(15 downto 0) := (others => '0');          -- number of bytes to transfer

    signal byte_count  : unsigned(15 downto 0) := (others => '0');          -- number of bytes transferred so far
    signal word_buf    : std_logic_vector(15 downto 0) := (others => '0');  -- buffer for the word to transfer

begin

    uart_controller: entity work.UART
        generic map (
            CLK_SPEED  => 50_000_000,     -- 50 MHz clock speed
            BAUD_RATE  => 38400           -- Baud rate for UART communication   -- (where two bytes is transferred in the time it takes to read/write a word in Spikeputor memory)
        )
        port map (
            CLK        => CLK,
            RST        => RST,
            RX_SERIAL  => UART_RXD,       -- Serial data input
            RX_DATA    => uart_rx_data,   -- Received byte output
            RX_READY   => uart_rx_rdy,    -- Strobed when a byte has been received
            TX_SERIAL  => UART_TXD,       -- Serial data output
            TX_DATA    => uart_tx_data,   -- Data to send through UART
            TX_LOAD    => uart_tx_load,   -- Strobe to send a byte
            TX_BUSY    => uart_tx_busy    -- Indicates if the transmitter is busy
        );



    -- flicker activity when the process is running, show completed when process is over and ready for next session
    ACTIVITY  <= '0' when (act_flasher < 25_000_000) else '1';
    COMPLETED <= '1' when (p_state = ACK_DONE OR p_state = WAIT_START) else '0';

    -- wire ADDR_OUT:
    ---    ADDR[21] is always 0
    ---    full sector address is 0 & ADDR[20:15] & 00000000000000
    ---    full address is 0 & sector address & (byte address/2)

    -- ADDR_OUT  <= ("0" & SECTOR_ADDR & "000000000000000") when (p_state = ERASE_FLASH OR p_state = WAIT_ERASE)
    --     else ("0" & SECTOR_ADDR & address);                                 -- set address to write to or sector to erase (when erase_flash was selected)
    ADDR_OUT  <= ("0" & address(20 downto 15) & "000000000000000") when (p_state = ERASE_FLASH OR p_state = WAIT_ERASE) AND address(20 downto 15) /= "000000"
            else "0000000111000000000000" when (p_state = ERASE_FLASH OR p_state = WAIT_ERASE) AND address(20 downto 15) = "000000"
            else ("0" & address);                                 -- set address to write to or sector to erase (when erase_flash was selected)

    -- wire DATA_OUT, WR_OUT and ERASE_OUT connections
    DATA_OUT  <= word_buf;                                                  -- set data to write
    WR_OUT    <= '1' when p_state = WRITE_FLASH else '0';                   -- strobe WR_OUT during the WRITE_FLASH state
    ERASE_OUT <= "10" when p_state = ERASE_FLASH else "00";                 -- strobe ERASE_OUT (to sector erase) during the ERASE_FLASH state

    --  State machine to implement transfer protocol
    process(CLK)
    begin
        if rising_edge(CLK) then
            TX_LOAD <= '0'; -- default TX_LOAD to '0'

            if RST = '1' then
                p_state <= WAIT_START;
                address <= (others => '0');
            else
                case (p_state) is

    --  WAIT_START: Wait for '*' or '?' to be recieved from UART
                    when WAIT_START =>                                      -- wait for RX_ready and rx_byte is '*'
                        if RX_READY = '1' then
                            if RX_DATA = C_STAR then
                                p_state <= ACK_UPLOAD;                      -- received '*', acknowledge by sending '!' and starting upload
                            elsif RX_DATA = C_QUES then
                                p_state <= ACK_ERASE;                       -- received '?', acknowledge by sending '!' and starting erase
                            end if;
                        end if;

    --  ACK_UPLOAD: Acknowledge the start of a new upload session with '!'
                    when ACK_UPLOAD =>
                        if TX_BUSY = '0' then
                            TX_DATA <=  C_BANG;
                            TX_LOAD <= '1';                                 -- strobe load signal (TX_DATA set above)
                            p_state <= HDR_0;                               -- start header read
                        end if;

    -- ACK_ERASE: Acknowledge the start of a new erase session with '!'
                    when ACK_ERASE =>
                        if TX_BUSY = '0' then
                            TX_DATA <= C_BANG;
                            TX_LOAD <= '1';                                 -- strobe load signal (TX_DATA set above)
                            p_state <= GET_SECTOR;                          -- start erase
                        end if;

    --  HDR_x: Read the 5 byte header (address, length) - address is byte address (22 bits), but low bit is ignored
                    when HDR_0 =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get high byte of address
                            address(20 downto 15) <= RX_DATA(5 downto 0);   -- store top 6 bits of byte address/2 = word address
                            p_state <= HDR_1;                               -- move to next header read state
                        end if;

                    when HDR_1 =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get next byte of address
                            address(14 downto 7) <= RX_DATA;                -- store next byte of byte address/2 = word address
                            p_state <= HDR_2;                               -- move to next header read state
                        end if;

                    when HDR_2 =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get low byte of address
                            address(6 downto 0) <= RX_DATA(7 downto 1);     -- store low byte of byte address/2 = word address
                            p_state <= HDR_3;                               -- move to next header read state
                        end if;

                    when HDR_3 =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get high byte of length of data
                            write_len(15 downto 8) <= unsigned(RX_DATA);    -- store high byte of length
                            p_state <= HDR_4;                               -- move to next header read state
                        end if;

                    when HDR_4 =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get low byte of length of data
                            write_len(7 downto 0) <= unsigned(RX_DATA);     -- store low byte of length
                            p_state <= LOAD_H;                              -- move to next state to load first word
                        end if;

    --  LOAD_x: read in two bytes of data to make the word to write to flash
                    when LOAD_H =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get high byte of word
                            word_buf(15 downto 8) <= RX_DATA;               -- store high byte of word
                            p_state  <= LOAD_L;                             -- move to next state to load low byte
                        end if;

                    when LOAD_L =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get low byte of word
                            word_buf(7 downto 0) <= RX_DATA;                -- store full word from byte_buf & low byte
                            p_state  <= WRITE_FLASH;                        -- move to next state to wait for flash to be ready to write
                        end if;

    -- WRITE_FLASH: write the word to flash at the current address
                    when WRITE_FLASH =>
                        if FLASH_RDY = '1' then
                            p_state   <= WAIT_FLASH;                        -- move to next state to wait for flash to finish writing
                        end if;

    -- WAIT_FLASH: wait for flash to be ready after it has written the word
                    when WAIT_FLASH =>
                        if FLASH_RDY = '1' then                             -- wait for flash idle
                            p_state <= NEXT_ADDRESS;                        -- move to next state to notify that flash has been written
                        end if;

    -- NEXT_ADDRESS: update address and byte counters, and check for end of data
                    when NEXT_ADDRESS =>
                        address     <= std_logic_vector(unsigned(address) + 1);     -- increment address by 1 (next word)
                        bytes_seen  <= bytes_seen + 2;                              -- increment byte counter by 2 (one word = 2 bytes)

                        if bytes_seen + 2 >= write_len then                 -- check if all data has been written
                            p_state <= ACK_DONE;                            -- if so, move to next state to acknowledge completion
                            bytes_seen <= (others => '0');                  -- and clear byte counter
                        else
                           p_state <= LOAD_H;                               -- otherwise, fetch next word
                    end if;

    -- GET_SECTOR: get sector to erase
                    when GET_SECTOR =>
                        if RX_READY = '1' then                              -- wait for RX_ready to get the 6 bit sector to erase
                            address(20 downto 15) <= RX_DATA(5 downto 0);   -- store top 6 bits of byte address/2 = word address
                            p_state <= ERASE_FLASH;                         -- move to next header read state
                        end if;

    -- ERASE_FLASH: send the command to erase the entire flash card
                    when ERASE_FLASH =>
                        if FLASH_RDY = '1' then
                            p_state <= WAIT_ERASE;                          -- move to the next state and wait for flash to finish erasing
                        end if;

    -- WAIT_ERASE: wait for flash to be ready after it erases the chip - increment counter so ACTIVITY light flashes at 1 Hz
                    when WAIT_ERASE =>
                        act_flasher <= act_flasher + 1;                -- increment activity counter, > 25_000_000 == ACTIVITY on

                        if act_flasher = 50_000_000 then
                            act_flasher <= 0;                               -- reset activity flasher at 50_000_000
                        end if;

                        if FLASH_RDY = '1' then                             -- wait for flash idle
                            act_flasher <= 0;                               -- reset the activity flasher counter
                            p_state <= ACK_DONE;                            -- move to next state to acknowledge completion
                        end if;

    --  ACK_DONE: send acknowledgement and reset state to wait for next upload
                    when ACK_DONE =>
                        if TX_BUSY = '0' then                               -- wait until UART is not busy to transmit
                            TX_DATA <=  C_STAR;
                            TX_LOAD <= '1';                                 -- strobe tx_load to transmit data
                            p_state <= WAIT_START;                          -- move to next state - ready for next session
                        end if;

                    when others =>
                        null;
                end case;
            end if;
        end if;
    end process;
end behavioral;